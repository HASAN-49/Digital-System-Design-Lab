module not_gate(x, y);
	input x;
	output y;
	not(y, x);
endmodule
